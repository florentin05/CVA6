/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module bootrom_64 (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic [63:0]  addr_i,
   output logic [63:0]  rdata_o
);
    localparam int RomSize = 918;

    const logic [RomSize-1:0][63:0] mem = {
        64'h00000000_00000000,
        64'h0a0d2165_6e6f6420,
        64'h00000000_00206567,
        64'h616d6920_746f6f62,
        64'h20676e69_79706f63,
        64'h00000000_00000009,
        64'h3a656d61_6e090a0d,
        64'h00093a73_65747562,
        64'h69727474_61090a0d,
        64'h00000009_3a61626c,
        64'h20747361_6c090a0d,
        64'h0000093a_61626c20,
        64'h74737269_66090a0d,
        64'h00000000_00000000,
        64'h09202020_20203a64,
        64'h69756720_6e6f6974,
        64'h69747261_70090a0d,
        64'h00000000_00000000,
        64'h093a6469_75672065,
        64'h70797420_6e6f6974,
        64'h69747261_70090a0d,
        64'h00000000_20797274,
        64'h6e65206e_6f697469,
        64'h74726170_20747067,
        64'h00000009_20203a73,
        64'h65697274_6e65206e,
        64'h6f697469_74726170,
        64'h20657a69_73090a0d,
        64'h00000009_3a736569,
        64'h72746e65_206e6f69,
        64'h74697472_61702072,
        64'h65626d75_6e090a0d,
        64'h00000009_2020203a,
        64'h61626c20_73656972,
        64'h746e6520_6e6f6974,
        64'h69747261_70090a0d,
        64'h00093a61_646c2070,
        64'h756b6361_62090a0d,
        64'h00000000_00000000,
        64'h093a6162_6c20746e,
        64'h65727275_63090a0d,
        64'h00000009_3a646576,
        64'h72657365_72090a0d,
        64'h00093a72_65646165,
        64'h685f6372_63090a0d,
        64'h00000000_00000909,
        64'h3a657a69_73090a0d,
        64'h00000009_3a6e6f69,
        64'h73697665_72090a0d,
        64'h0000093a_65727574,
        64'h616e6769_73090a0d,
        64'h00000000_003a7265,
        64'h64616568_20656c62,
        64'h6174206e_6f697469,
        64'h74726170_20747067,
        64'h0000203a_65756c61,
        64'h76206e72_75746572,
        64'h2079706f_63206473,
        64'h00000000_0000000a,
        64'h0d216465_6c696166,
        64'h20647261_63204453,
        64'h00000000_0000000a,
        64'h0d216465_7a696c61,
        64'h6974696e_69206473,
        64'h00000000_0a0d676e,
        64'h69746978_65202e2e,
        64'h2e647320_657a696c,
        64'h61697469_6e692074,
        64'h6f6e2064_6c756f63,
        64'h00000000_0000002e,
        64'h00000000_0000000a,
        64'h0d6b636f_6c622044,
        64'h53206461_65722074,
        64'h6f6e2064_6c756f63,
        64'h0000000a_0d202e2e,
        64'h2e445320_676e697a,
        64'h696c6169_74696e69,
        64'h00000031_34646d63,
        64'h00000035_35646d63,
        64'h00000000_30646d63,
        64'h00000020_3a206573,
        64'h6e6f7073_65720920,
        64'h00000000_0020646e,
        64'h616d6d6f_63204453,
        64'h00000000_203f3f79,
        64'h74706d65_20746f6e,
        64'h206f6669_66207872,
        64'h00000000_00000a0d,
        64'h2164657a_696c6169,
        64'h74696e69_20495053,
        64'h00000000_00007830,
        64'h203a7375_74617473,
        64'h00000000_00000a0d,
        64'h49505320_74696e69,
        64'h00000000_000a0d33,
        64'h3230322c_49534149,
        64'h00000000_00000000,
        64'h0a0d6965_72646e41,
        64'h204e4154_53202e67,
        64'h6e49202e_7244202e,
        64'h666f7250_203a726f,
        64'h74616d75_72646e49,
        64'h00000000_0000000a,
        64'h0d6e6974_6e65726f,
        64'h6c462045_494c4920,
        64'h3a746e65_64757453,
        64'h00000000_000a0d56,
        64'h2d435349_5220696e,
        64'h75697463_75727473,
        64'h6e692065_64206c75,
        64'h74657320_646e617a,
        64'h696c6974_7520436f,
        64'h53206975_6e752061,
        64'h65726174_6365696f,
        64'h7250203a_74636569,
        64'h6f727020_616d6554,
        64'h00000000_0000000a,
        64'h0d414d4f_4c504944,
        64'h20746365_696f7250,
        64'h00000000_00000032,
        64'h2d746c75_61666564,
        64'h2d697274_2c786e6c,
        64'h7800746c_75616665,
        64'h642d6972_742c786e,
        64'h6c78006c_6175642d,
        64'h73692c78_6e6c7800,
        64'h746e6573_6572702d,
        64'h74707572_7265746e,
        64'h692c786e_6c780068,
        64'h74646977_2d326f69,
        64'h70672c78_6e6c7800,
        64'h68746469_772d6f69,
        64'h70672c78_6e6c7800,
        64'h322d746c_75616665,
        64'h642d7475_6f642c78,
        64'h6e6c7800_746c7561,
        64'h6665642d_74756f64,
        64'h2c786e6c_7800322d,
        64'h73747570_6e692d6c,
        64'h6c612c78_6e6c7800,
        64'h73747570_6e692d6c,
        64'h6c612c78_6e6c7800,
        64'h72656c6c_6f72746e,
        64'h6f632d6f_69706700,
        64'h736c6c65_632d6f69,
        64'h70672300_73736572,
        64'h6464612d_63616d2d,
        64'h6c61636f_6c007077,
        64'h2d656c62_61736964,
        64'h00736567_6e61722d,
        64'h65676174_6c6f7600,
        64'h79636e65_75716572,
        64'h662d7861_6d2d6970,
        64'h73006f69_7461722d,
        64'h6b63732c_786e6c78,
        64'h00737469_622d7265,
        64'h66736e61_72742d6d,
        64'h756e2c78_6e6c7800,
        64'h73746962_2d73732d,
        64'h6d756e2c_786e6c78,
        64'h00747369_78652d6f,
        64'h6669662c_786e6c78,
        64'h00796c69_6d61662c,
        64'h786e6c78_00687464,
        64'h69772d6f_692d6765,
        64'h72007466_6968732d,
        64'h67657200_73747075,
        64'h72726574_6e690074,
        64'h6e657261_702d7470,
        64'h75727265_746e6900,
        64'h64656570_732d746e,
        64'h65727275_63007665,
        64'h646e2c76_63736972,
        64'h00797469_726f6972,
        64'h702d7861_6d2c7663,
        64'h73697200_73656d61,
        64'h6e2d6765_72006465,
        64'h646e6574_78652d73,
        64'h74707572_7265746e,
        64'h69007365_676e6172,
        64'h00646564_6e657073,
        64'h75732d65_74617473,
        64'h2d6e6961_74657200,
        64'h72656767_6972742d,
        64'h746c7561_6665642c,
        64'h78756e69_6c00736f,
        64'h69706700_656c646e,
        64'h61687000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h00736c6c_65632d74,
        64'h70757272_65746e69,
        64'h23007469_6c70732d,
        64'h626c7400_65707974,
        64'h2d756d6d_00617369,
        64'h2c766373_69720073,
        64'h75746174_73006765,
        64'h72006570_79745f65,
        64'h63697665_64007963,
        64'h6e657571_6572662d,
        64'h6b636f6c_63007963,
        64'h6e657571_6572662d,
        64'h65736162_656d6974,
        64'h00687461_702d7475,
        64'h6f647473_006c6564,
        64'h6f6d0065_6c626974,
        64'h61706d6f_6300736c,
        64'h6c65632d_657a6973,
        64'h2300736c_6c65632d,
        64'h73736572_64646123,
        64'h09000000_02000000,
        64'h02000000_02000000,
        64'h01000000_b5000000,
        64'h04000000_03000000,
        64'hffffffff_bf020000,
        64'h04000000_03000000,
        64'hffffffff_ae020000,
        64'h04000000_03000000,
        64'h01000000_a1020000,
        64'h04000000_03000000,
        64'h00000000_8a020000,
        64'h04000000_03000000,
        64'h08000000_79020000,
        64'h04000000_03000000,
        64'h08000000_69020000,
        64'h04000000_03000000,
        64'h00000000_55020000,
        64'h04000000_03000000,
        64'h00000000_43020000,
        64'h04000000_03000000,
        64'h00000000_31020000,
        64'h04000000_03000000,
        64'h00000000_21020000,
        64'h04000000_03000000,
        64'h00000100_00000000,
        64'h00000040_00000000,
        64'h67000000_10000000,
        64'h03000000_11020000,
        64'h00000000_03000000,
        64'h00000000_612e3030,
        64'h2e312d6f_6970672d,
        64'h7370782c_786e6c78,
        64'h1b000000_15000000,
        64'h03000000_02000000,
        64'h05020000_04000000,
        64'h03000000_00000030,
        64'h30303030_30303440,
        64'h6f697067_01000000,
        64'h02000000_00800000,
        64'h00000000_00000030,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h00007fe3_023e1800,
        64'hf3010000_06000000,
        64'h03000000_00000000,
        64'h03000000_52010000,
        64'h08000000_03000000,
        64'h03000000_41010000,
        64'h04000000_03000000,
        64'h006b726f_7774656e,
        64'h5b000000_08000000,
        64'h03000000_00687465,
        64'h2d637369_72776f6c,
        64'h1b000000_0c000000,
        64'h03000000_00000000,
        64'h30303030_30303033,
        64'h40687465_2d637369,
        64'h72776f6c_01000000,
        64'h02000000_02000000,
        64'he8010000_00000000,
        64'h03000000_e40c0000,
        64'he40c0000_d9010000,
        64'h08000000_03000000,
        64'h20bcbe00_c7010000,
        64'h04000000_03000000,
        64'h00000000_67000000,
        64'h04000000_03000000,
        64'h00000000_746f6c73,
        64'h2d697073_2d636d6d,
        64'h1b000000_0d000000,
        64'h03000000_00000030,
        64'h40636d6d_01000000,
        64'h04000000_b8010000,
        64'h04000000_03000000,
        64'h08000000_a1010000,
        64'h04000000_03000000,
        64'h01000000_90010000,
        64'h04000000_03000000,
        64'h01000000_80010000,
        64'h04000000_03000000,
        64'h00377865_746e696b,
        64'h74010000_08000000,
        64'h03000000_00100000,
        64'h00000000_00000020,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h02000000_02000000,
        64'h52010000_08000000,
        64'h03000000_03000000,
        64'h41010000_04000000,
        64'h03000000_00000000,
        64'h0f000000_04000000,
        64'h03000000_01000000,
        64'h00000000_04000000,
        64'h03000000_00612e30,
        64'h302e322d_6970732d,
        64'h7370782c_786e6c78,
        64'h00622e30_302e322d,
        64'h6970732d_7370782c,
        64'h786e6c78_1b000000,
        64'h28000000_03000000,
        64'h00000000_30303030,
        64'h30303032_40697073,
        64'h2d737078_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_0b010000,
        64'h08000000_03000000,
        64'h03000000_41010000,
        64'h04000000_03000000,
        64'h00100000_00000000,
        64'h00000018_00000000,
        64'h67000000_10000000,
        64'h03000000_07000000,
        64'h06000000_05000000,
        64'h04000000_52010000,
        64'h10000000_03000000,
        64'h00007265_6d69745f,
        64'h6270612c_706c7570,
        64'h1b000000_0f000000,
        64'h03000000_00003030,
        64'h30303030_38314072,
        64'h656d6974_01000000,
        64'h02000000_04000000,
        64'h67010000_04000000,
        64'h03000000_02000000,
        64'h5d010000_04000000,
        64'h03000000_01000000,
        64'h52010000_04000000,
        64'h03000000_03000000,
        64'h41010000_04000000,
        64'h03000000_00c20100,
        64'h33010000_04000000,
        64'h03000000_80f0fa02,
        64'h4b000000_04000000,
        64'h03000000_00100000,
        64'h00000000_00000010,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h00000000_61303535,
        64'h3631736e_1b000000,
        64'h09000000_03000000,
        64'h00000030_30303030,
        64'h30303140_74726175,
        64'h01000000_02000000,
        64'h03000000_b5000000,
        64'h04000000_03000000,
        64'h1e000000_28010000,
        64'h04000000_03000000,
        64'h07000000_15010000,
        64'h04000000_03000000,
        64'h00000004_00000000,
        64'h0000000c_00000000,
        64'h67000000_10000000,
        64'h03000000_09000000,
        64'h02000000_0b000000,
        64'h02000000_f7000000,
        64'h10000000_03000000,
        64'ha0000000_00000000,
        64'h03000000_00306369,
        64'h6c702c76_63736972,
        64'h1b000000_0c000000,
        64'h03000000_01000000,
        64'h8f000000_04000000,
        64'h03000000_00000000,
        64'h00000000_04000000,
        64'h03000000_00000000,
        64'h30303030_30306340,
        64'h72656c6c_6f72746e,
        64'h6f632d74_70757272,
        64'h65746e69_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_0b010000,
        64'h08000000_03000000,
        64'h00000c00_00000000,
        64'h00000002_00000000,
        64'h67000000_10000000,
        64'h03000000_07000000,
        64'h02000000_03000000,
        64'h02000000_f7000000,
        64'h10000000_03000000,
        64'h00000000_30746e69,
        64'h6c632c76_63736972,
        64'h1b000000_0d000000,
        64'h03000000_00000030,
        64'h30303030_30324074,
        64'h6e696c63_01000000,
        64'hf0000000_00000000,
        64'h03000000_00007375,
        64'h622d656c_706d6973,
        64'h00636f73_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h1f000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00636f73_01000000,
        64'h02000000_02000000,
        64'hd9000000_00000000,
        64'h03000000_00000074,
        64'h61656274_72616568,
        64'hc3000000_0a000000,
        64'h03000000_00000000,
        64'h01000000_01000000,
        64'hbd000000_0c000000,
        64'h03000000_00000064,
        64'h656c2d74_61656274,
        64'h72616568_01000000,
        64'h00000073_64656c2d,
        64'h6f697067_1b000000,
        64'h0a000000_03000000,
        64'h00000000_7364656c,
        64'h01000000_02000000,
        64'h00000040_00000000,
        64'h00000080_00000000,
        64'h67000000_10000000,
        64'h03000000_00007972,
        64'h6f6d656d_5b000000,
        64'h07000000_03000000,
        64'h00303030_30303030,
        64'h38407972_6f6d656d,
        64'h01000000_02000000,
        64'h02000000_02000000,
        64'h02000000_b5000000,
        64'h04000000_03000000,
        64'h00006374_6e692d75,
        64'h70632c76_63736972,
        64'h1b000000_0f000000,
        64'h03000000_a0000000,
        64'h00000000_03000000,
        64'h01000000_8f000000,
        64'h04000000_03000000,
        64'h00000000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h01000000_85000000,
        64'h00000000_03000000,
        64'h00003933_76732c76,
        64'h63736972_7c000000,
        64'h0b000000_03000000,
        64'h00006364_66616d69,
        64'h34367672_72000000,
        64'h0b000000_03000000,
        64'h00000076_63736972,
        64'h00656e61_69726120,
        64'h2c687465_1b000000,
        64'h12000000_03000000,
        64'h00000000_79616b6f,
        64'h6b000000_05000000,
        64'h03000000_00000000,
        64'h67000000_04000000,
        64'h03000000_00757063,
        64'h5b000000_04000000,
        64'h03000000_80f0fa02,
        64'h4b000000_04000000,
        64'h03000000_00000030,
        64'h40757063_01000000,
        64'h40787d01_38000000,
        64'h04000000_03000000,
        64'h00000000_0f000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00000000_73757063,
        64'h01000000_02000000,
        64'h00000030_30323531,
        64'h313a3030_30303030,
        64'h30314074_7261752f,
        64'h636f732f_2c000000,
        64'h1a000000_03000000,
        64'h00006e65_736f6863,
        64'h01000000_00657261,
        64'h622d656e_61697261,
        64'h2c687465_26000000,
        64'h10000000_03000000,
        64'h00766564_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h14000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00000000_01000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'he8080000_d2020000,
        64'h00000000_10000000,
        64'h11000000_28000000,
        64'h20090000_38000000,
        64'hf20b0000_edfe0dd0,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h46454443_42413938,
        64'h37363534_33323130,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'hbfe1c63e_37fd47b2,
        64'hbfc90091_05a3ffe1,
        64'h0ff7f793_00b14783,
        64'h00f105a3_838500b1,
        64'h478300f0_4f632781,
        64'h47b2c622_f73ff0ef,
        64'h40000537_00b14583,
        64'h54fdf8df_f0ef5a04,
        64'h0413e68f_f0ef0026,
        64'h2437eb25_05130000,
        64'h1517e78f_f0efe8e5,
        64'h05130000_1517e84f,
        64'hf0efe7a5_05130000,
        64'h1517e90f_f0efe365,
        64'h05130000_1517e9cf,
        64'hf0efe2a5_05130000,
        64'h1517e64f_f0efec26,
        64'hf02200f1_05a3f406,
        64'h08050513_20058593,
        64'h57fd7179_02faf537,
        64'h65f18082_00e78623,
        64'h477d0007_82234000,
        64'h07b78082_00054503,
        64'h808200b5_0023bbb9,
        64'hee6ff0ef_21c50513,
        64'h00001517_bbc1f765,
        64'h05130000_1517f7ef,
        64'hf0ef8526_f02ff0ef,
        64'h07850513_00001517,
        64'hf0eff0ef_06c50513,
        64'h00001517_bbe5f9e5,
        64'h05130000_1517fa6f,
        64'hf0ef8526_f2aff0ef,
        64'h0a050513_00001517,
        64'hf36ff0ef_09450513,
        64'h00001517_c92984aa,
        64'hc3dff0ef_9e0d2605,
        64'h855a020a_a583028a,
        64'hb603f58f_f0ef2765,
        64'h05130000_1517f374,
        64'h9de30809_09130809,
        64'h8993f70f_f0ef2485,
        64'hff850513_00001517,
        64'hff499be3_847ff0ef,
        64'h0a05000a_4503f8cf,
        64'hf0ef29a5_05130000,
        64'h151781bf_f0ef0109,
        64'h3503fa0f_f0ef29e5,
        64'h05130000_151782ff,
        64'hf0ef0089_3503fb4f,
        64'hf0ef2a25_05130000,
        64'h1517843f_f0effb89,
        64'h8a130009_3503fccf,
        64'hf0ef2aa5_05130000,
        64'h1517ff2a_1be38a1f,
        64'hf0ef0a05_000a4503,
        64'hf9098a13_feaff0ef,
        64'h2a850513_00001517,
        64'hff8a19e3_8bfff0ef,
        64'h0a050007_c503014c,
        64'h87b34a01_80bff0ef,
        64'hf8098c93_2ac50513,
        64'h00001517_8dfff0ef,
        64'h0ff4f513_823ff0ef,
        64'h2a850513_00001517,
        64'h4b914c41_10051e63,
        64'h02010913_08010993,
        64'h84aa8a8a_d39ff0ef,
        64'h850a4605_71010489,
        64'h2583851f_f0ef0d65,
        64'h05130000_151789ff,
        64'hf0ef4556_863ff0ef,
        64'h2c850513_00001517,
        64'h8b1ff0ef_4546875f,
        64'hf0ef2ba5_05130000,
        64'h1517903f_f0ef6526,
        64'h887ff0ef_2ac50513,
        64'h00001517_915ff0ef,
        64'h7502899f_f0ef2ae5,
        64'h05130000_1517927f,
        64'hf0ef6562_8abff0ef,
        64'h2a850513_00001517,
        64'h8f9ff0ef_45528bdf,
        64'hf0ef2aa5_05130000,
        64'h151790bf_f0ef4542,
        64'h8cfff0ef_2ac50513,
        64'h00001517_91dff0ef,
        64'h45328e1f_f0ef2ae5,
        64'h05130000_151792ff,
        64'hf0ef4522_8f3ff0ef,
        64'h2b050513_00001517,
        64'h981ff0ef_6502905f,
        64'hf0ef2b25_05130000,
        64'h1517911f_f0ef29e5,
        64'h05130000_1517bf59,
        64'h54f9921f_f0ef1a65,
        64'h05130000_15179aff,
        64'hf0ef8526_933ff0ef,
        64'h2a850513_00001517,
        64'h93fff0ef_29c50513,
        64'h00001517_c90584aa,
        64'h890ae47f_f0ef850a,
        64'h45854605_710195df,
        64'hf0ef2a25_05130000,
        64'h15178082_61256ca2,
        64'h6c426be2_7b027aa2,
        64'h7a4279e2_690664a6,
        64'h64468526_60e6fa04,
        64'h011354fd_98bff0ef,
        64'h2a850513_00001517,
        64'hc905df3f_f0ef8b2a,
        64'h1080e466_e862ec5e,
        64'hf456f852_fc4ee0ca,
        64'he4a6ec86_f05ae8a2,
        64'h711db765_54798082,
        64'h61696baa_6b4a6aea,
        64'h7a0a79aa_794a74ea,
        64'h640e60ae_8522547d,
        64'h9d7ff0ef_2cc50513,
        64'h00001517_c61ff0ef,
        64'hc65ff0ef_c69ff0ef,
        64'hc6dff0ef_c71ff0ef,
        64'hc75ff0ef_c79ff0ef,
        64'hc7dff0ef_a805c83f,
        64'hf0efc8df_f0ef4531,
        64'h45814605_4401f930,
        64'h46e32004_849319fd,
        64'ha1fff0ef_33450513,
        64'h00001517_e7990369,
        64'he7b30689_1c639041,
        64'h29011442_8c49cbbf,
        64'hf0ef9041_03051413,
        64'h0085151b_cc9ff0ef,
        64'hfc941ae3_04040413,
        64'hff7a17e3_892af15f,
        64'hf0ef0a05_854a0007,
        64'hc5830144_07b30400,
        64'h0b934a01_c6dff0ef,
        64'h850a0400_05938622,
        64'h4901ff55_1ee3d03f,
        64'hf0efe004_84133e80,
        64'h0b130fe0_0a93e951,
        64'h20048493_d1fff0ef,
        64'h454985a2_0ff67613,
        64'h00166613_0015161b,
        64'hf4dff0ef_0ff47593,
        64'hf55ff0ef_0ff5f593,
        64'h0084559b_f61ff0ef,
        64'h0ff5f593_0104559b,
        64'hf6dff0ef_45010184,
        64'h559bfee7_9be30785,
        64'h00c68023_00f106b3,
        64'h08000713_567d4781,
        64'h0209d993_842e84aa,
        64'he55ee95a_ed56f152,
        64'hf94ae586_fd26e1a2,
        64'h02061993_f54e7155,
        64'h80829141_15428d3d,
        64'h8ff90057_979b1701,
        64'h67090107_d79b0105,
        64'h179b4105_551b0105,
        64'h151b8d2d_00c59513,
        64'h8da9893d_0045d51b,
        64'h8da99141_15428d5d,
        64'h05220085_579b8082,
        64'h07f57513_8d2d0045,
        64'h15938d2d_8d3d0045,
        64'hd51b0075_d79b8de9,
        64'h80820141_853e6402,
        64'h60a257f5_e1114781,
        64'hf89ff0ef_c51157f9,
        64'hefbff0ef_c91157fd,
        64'heb7ff0ef_fc6de0bf,
        64'hf0ef347d_4429b95f,
        64'hf0ef4725_05130000,
        64'h1517c8ff_f0efe022,
        64'he4061141_80826105,
        64'h00153513_64a26442,
        64'h60e20004_051bfc94,
        64'h0ce3e3ff_f0efeb5f,
        64'hf0ef49a5_05130000,
        64'h151785aa_842ae59f,
        64'hf0ef0290_05134000,
        64'h05b70770_0613fbdf,
        64'hf0ef4485_e822ec06,
        64'he4261101_80820141,
        64'h00153513_157d6402,
        64'h60a20004_051bef5f,
        64'hf0ef4d45_051385a2,
        64'h00001517_e91ff0ef,
        64'h842ae9df_f0efe022,
        64'he4060370_05134581,
        64'h06500613_11418082,
        64'h61056902_64a26442,
        64'h60e20015_3513f565,
        64'h05130004_051b0124,
        64'h986388bd_00f91b63,
        64'h45014785_ed1ff0ef,
        64'hed5ff0ef_842aedbf,
        64'hf0ef84aa_ee1ff0ef,
        64'hee5ff0ef_ee9ff0ef,
        64'h892aef5f_f0efe04a,
        64'he426e822_ec064521,
        64'h1aa00593_08700613,
        64'h1101bfcd_45018082,
        64'h61056902_64a26442,
        64'h60e24505_f8bff0ef,
        64'h45855625_05130000,
        64'h1517fe99_15e3c00d,
        64'hf2dff0ef_892a347d,
        64'hf3bff0ef_45014581,
        64'h09500613_44857104,
        64'h0413e04a_ec06e426,
        64'h6409e822_1101b9c9,
        64'h610555a5_05130000,
        64'h151760e2_6442da9f,
        64'hf0ef852e_65a2cedf,
        64'hf0ef5a25_05130000,
        64'h1517cf9f_f0ef8522,
        64'hcffff0ef_e42eec06,
        64'h5a850513_00001517,
        64'h842ae822_11018082,
        64'h614564e2_740270a2,
        64'hf47d147d_0007d463,
        64'h4187d79b_0185179b,
        64'hfadff0ef_eb7ff0ef,
        64'h85320640_04136622,
        64'hec3ff0ef_0ff47513,
        64'hecbff0ef_0ff57513,
        64'h0084551b_ed7ff0ef,
        64'h0ff57513_0104551b,
        64'hee3ff0ef_0184551b,
        64'heebff0ef_0404e513,
        64'hfedff0ef_84aa842e,
        64'hec26f022_e432f406,
        64'h7179b709_0ff00513,
        64'h8082557d_b7d900d7,
        64'h00230785_00f60733,
        64'h06c82683_ff698b05,
        64'h5178b77d_d6b80785,
        64'h00074703_00f50733,
        64'h80824501_d3b84719,
        64'hdbb8577d_200007b7,
        64'h02b6e163_0007869b,
        64'h20000837_20000537,
        64'hfff58b85_537c2000,
        64'h0737d3b8_200007b7,
        64'h10600713_fff537fd,
        64'h00010320_079304b7,
        64'h61630007_871b4781,
        64'h200006b7_dbb85779,
        64'h200007b7_06b7ee63,
        64'h10000793_80826105,
        64'h64a2d3b8_4719dbb8,
        64'h644260e2_0ff47513,
        64'h577d2000_07b7e25f,
        64'hf0ef6aa5_05130000,
        64'h1517eb3f_f0ef9101,
        64'h15024088_e3bff0ef,
        64'h6c850513_00001517,
        64'he3958b85_240153fc,
        64'h57e0ff65_8b050647,
        64'h849353f8_d3b81060,
        64'h07132000_07b7fff5,
        64'h37fd0001_06400793,
        64'hd7a8dbb8_5779e426,
        64'he822ec06_200007b7,
        64'h1101bdbd_61056f65,
        64'h05130000_151764a2,
        64'h60e26442_d03c4799,
        64'he97ff0ef_71c50513,
        64'h00001517_f25ff0ef,
        64'h91010204_95132481,
        64'heafff0ef_71450513,
        64'h00001517_5064d03c,
        64'h16600793_ec3ff0ef,
        64'h74850513_00001517,
        64'hf51ff0ef_91010204,
        64'h95132481_edbff0ef,
        64'h74050513_00001517,
        64'h5064d03c_10400793,
        64'h20000437_fff537fd,
        64'h000147a9_c3b84729,
        64'h200007b7_f03ff0ef,
        64'he426e822_ec067605,
        64'h05131101_00001517,
        64'h80822501_41088082,
        64'hc10c8082_610560e2,
        64'hecfff0ef_00914503,
        64'hed7ff0ef_00814503,
        64'hf55ff0ef_ec06002c,
        64'h11018082_61456942,
        64'h64e27402_70a2fe94,
        64'h10e3ef9f_f0ef0091,
        64'h4503f01f_f0ef3461,
        64'h00814503_f81ff0ef,
        64'h0ff57513_002c0089,
        64'h553354e1_03800413,
        64'h892af406_e84aec26,
        64'hf0227179_80826145,
        64'h694264e2_740270a2,
        64'hfe9410e3_f3bff0ef,
        64'h00914503_f43ff0ef,
        64'h34610081_4503fc3f,
        64'hf0ef0ff5_7513002c,
        64'h0089553b_54e14461,
        64'h892af406_e84aec26,
        64'hf0227179_808200f5,
        64'h80230007_c78300e5,
        64'h80a397aa_81110007,
        64'h4703973e_00f57713,
        64'ha7078793_00001797,
        64'hb7f50405_f93ff0ef,
        64'h80820141_640260a2,
        64'he5090004_4503842a,
        64'he406e022_11418082,
        64'h00e78823_02000713,
        64'h00e78423_fc700713,
        64'h00e78623_470d00a7,
        64'h82230ff5_751300e7,
        64'h80230085_551b0ff5,
        64'h771300e7_8623f800,
        64'h07130007_82231000,
        64'h07b702b5_553b0045,
        64'h959b8082_00a70023,
        64'hdfe50207_f7930147,
        64'h47831000_07378082,
        64'h02057513_0147c503,
        64'h100007b7_80820005,
        64'h45038082_00b50023,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00048067_01f49493,
        64'h0010049b_c8458593,
        64'h00001597_f1402573,
        64'hff24c6e3_4009091b,
        64'h02000937_00448493,
        64'hfe091ee3_0004a903,
        64'h00092023_00990933,
        64'h00291913_f1402973,
        64'h020004b7_fe090ae3,
        64'h00897913_34402973,
        64'h10500073_ff24c6e3,
        64'h4009091b_02000937,
        64'h00448493_0124a023,
        64'h00100913_020004b7,
        64'h293000ef_01a11113,
        64'h0210011b_03249663,
        64'hf1402973_00000493,
        64'h30491073_00800913
    };

    logic [$clog2(RomSize)-1:0] addr_q;

    always_ff @(posedge clk_i) begin
        if (req_i) begin
            addr_q <= addr_i[$clog2(RomSize)-1+3:3];
        end
    end

    // this prevents spurious Xes from propagating into
    // the speculative fetch stage of the core
    assign rdata_o = (addr_q < RomSize) ? mem[addr_q] : '0;
endmodule
