/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module bootrom_64 (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic [63:0]  addr_i,
   output logic [63:0]  rdata_o
);
    localparam int RomSize = 1081;

    const logic [RomSize-1:0][63:0] mem = {
        64'hfffefdfc_fbfaf9f8,
        64'h00000000_00000000,
        64'h0a0d2165_6e6f6420,
        64'h00000000_00206567,
        64'h616d6920_746f6f62,
        64'h20676e69_79706f63,
        64'h00000000_00000009,
        64'h3a656d61_6e090a0d,
        64'h00093a73_65747562,
        64'h69727474_61090a0d,
        64'h00000009_3a61626c,
        64'h20747361_6c090a0d,
        64'h0000093a_61626c20,
        64'h74737269_66090a0d,
        64'h00000000_00000000,
        64'h09202020_20203a64,
        64'h69756720_6e6f6974,
        64'h69747261_70090a0d,
        64'h00000000_00000000,
        64'h093a6469_75672065,
        64'h70797420_6e6f6974,
        64'h69747261_70090a0d,
        64'h00000000_20797274,
        64'h6e65206e_6f697469,
        64'h74726170_20747067,
        64'h00000009_20203a73,
        64'h65697274_6e65206e,
        64'h6f697469_74726170,
        64'h20657a69_73090a0d,
        64'h00000009_3a736569,
        64'h72746e65_206e6f69,
        64'h74697472_61702072,
        64'h65626d75_6e090a0d,
        64'h00000009_2020203a,
        64'h61626c20_73656972,
        64'h746e6520_6e6f6974,
        64'h69747261_70090a0d,
        64'h00093a61_646c2070,
        64'h756b6361_62090a0d,
        64'h00000000_00000000,
        64'h093a6162_6c20746e,
        64'h65727275_63090a0d,
        64'h00000009_3a646576,
        64'h72657365_72090a0d,
        64'h00093a72_65646165,
        64'h685f6372_63090a0d,
        64'h00000000_00000909,
        64'h3a657a69_73090a0d,
        64'h00000009_3a6e6f69,
        64'h73697665_72090a0d,
        64'h0000093a_65727574,
        64'h616e6769_73090a0d,
        64'h00000000_003a7265,
        64'h64616568_20656c62,
        64'h6174206e_6f697469,
        64'h74726170_20747067,
        64'h0000203a_65756c61,
        64'h76206e72_75746572,
        64'h2079706f_63206473,
        64'h00000000_0000000a,
        64'h0d216465_6c696166,
        64'h20647261_63204453,
        64'h00000000_0000000a,
        64'h0d216465_7a696c61,
        64'h6974696e_69206473,
        64'h00000000_0a0d676e,
        64'h69746978_65202e2e,
        64'h2e647320_657a696c,
        64'h61697469_6e692074,
        64'h6f6e2064_6c756f63,
        64'h00000000_0000002e,
        64'h00000000_0000000a,
        64'h0d6b636f_6c622044,
        64'h53206461_65722074,
        64'h6f6e2064_6c756f63,
        64'h0000000a_0d202e2e,
        64'h2e445320_676e697a,
        64'h696c6169_74696e69,
        64'h00000031_34646d63,
        64'h00000035_35646d63,
        64'h00000000_30646d63,
        64'h00000020_3a206573,
        64'h6e6f7073_65720920,
        64'h00000000_0020646e,
        64'h616d6d6f_63204453,
        64'h00000000_203f3f79,
        64'h74706d65_20746f6e,
        64'h206f6669_66207872,
        64'h00000000_00000a0d,
        64'h2164657a_696c6169,
        64'h74696e69_20495053,
        64'h00000000_00007830,
        64'h203a7375_74617473,
        64'h00000000_00000a0d,
        64'h49505320_74696e69,
        64'h0000003a_4d415220,
        64'h6e696420_69726974,
        64'h69632030_30303030,
        64'h31207470_20696c63,
        64'h6963202e_724e0a0d,
        64'h0000003a_4d415220,
        64'h6e692069_72656972,
        64'h63732030_30303030,
        64'h31207470_20696c63,
        64'h6963202e_724e0a0d,
        64'h00000000_3a4d4152,
        64'h206e6964_20697269,
        64'h74696320_30303030,
        64'h31207470_20696c63,
        64'h6963202e_724e0a0d,
        64'h00000000_3a4d4152,
        64'h206e6920_69726569,
        64'h72637320_30303030,
        64'h31207470_20696c63,
        64'h6963202e_724e0a0d,
        64'h00000000_00003a4d,
        64'h4152206e_69642069,
        64'h72697469_63203030,
        64'h31207470_20696c63,
        64'h6963202e_724e0a0d,
        64'h00000000_00003a4d,
        64'h4152206e_69206972,
        64'h65697263_73203030,
        64'h31207470_20696c63,
        64'h6963202e_724e0a0d,
        64'h000a0d20_65697469,
        64'h72617061_20616d69,
        64'h7270203a_454e5549,
        64'h54435552_54534e49,
        64'h00000a0d_20623878,
        64'h616d203a_454e5549,
        64'h54435552_54534e49,
        64'h00000000_00000000,
        64'h203a696c_63696320,
        64'h74726f70_61520a0d,
        64'h00000000_0000203a,
        64'h656e7569_74637572,
        64'h74736e69_20696c63,
        64'h6963202e_724e0a0d,
        64'h00000000_00203a43,
        64'h20646f63_20696c63,
        64'h6963202e_724e0a0d,
        64'h00000000_00000000,
        64'h203a656e_75697463,
        64'h75727473_6e692073,
        64'h6e757073_61520a0d,
        64'h00203a43_20646f63,
        64'h20736e75_70736152,
        64'h00000000_000a0d20,
        64'h73656e6f_5f746e75,
        64'h6f63203a_454e5549,
        64'h54435552_54534e49,
        64'h00000a0d_21646c72,
        64'h6f57206f_6c6c6548,
        64'h00000000_00000032,
        64'h2d746c75_61666564,
        64'h2d697274_2c786e6c,
        64'h7800746c_75616665,
        64'h642d6972_742c786e,
        64'h6c78006c_6175642d,
        64'h73692c78_6e6c7800,
        64'h746e6573_6572702d,
        64'h74707572_7265746e,
        64'h692c786e_6c780068,
        64'h74646977_2d326f69,
        64'h70672c78_6e6c7800,
        64'h68746469_772d6f69,
        64'h70672c78_6e6c7800,
        64'h322d746c_75616665,
        64'h642d7475_6f642c78,
        64'h6e6c7800_746c7561,
        64'h6665642d_74756f64,
        64'h2c786e6c_7800322d,
        64'h73747570_6e692d6c,
        64'h6c612c78_6e6c7800,
        64'h73747570_6e692d6c,
        64'h6c612c78_6e6c7800,
        64'h72656c6c_6f72746e,
        64'h6f632d6f_69706700,
        64'h736c6c65_632d6f69,
        64'h70672300_73736572,
        64'h6464612d_63616d2d,
        64'h6c61636f_6c007077,
        64'h2d656c62_61736964,
        64'h00736567_6e61722d,
        64'h65676174_6c6f7600,
        64'h79636e65_75716572,
        64'h662d7861_6d2d6970,
        64'h73006f69_7461722d,
        64'h6b63732c_786e6c78,
        64'h00737469_622d7265,
        64'h66736e61_72742d6d,
        64'h756e2c78_6e6c7800,
        64'h73746962_2d73732d,
        64'h6d756e2c_786e6c78,
        64'h00747369_78652d6f,
        64'h6669662c_786e6c78,
        64'h00796c69_6d61662c,
        64'h786e6c78_00687464,
        64'h69772d6f_692d6765,
        64'h72007466_6968732d,
        64'h67657200_73747075,
        64'h72726574_6e690074,
        64'h6e657261_702d7470,
        64'h75727265_746e6900,
        64'h64656570_732d746e,
        64'h65727275_63007665,
        64'h646e2c76_63736972,
        64'h00797469_726f6972,
        64'h702d7861_6d2c7663,
        64'h73697200_73656d61,
        64'h6e2d6765_72006465,
        64'h646e6574_78652d73,
        64'h74707572_7265746e,
        64'h69007365_676e6172,
        64'h00646564_6e657073,
        64'h75732d65_74617473,
        64'h2d6e6961_74657200,
        64'h72656767_6972742d,
        64'h746c7561_6665642c,
        64'h78756e69_6c00736f,
        64'h69706700_656c646e,
        64'h61687000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h00736c6c_65632d74,
        64'h70757272_65746e69,
        64'h23007469_6c70732d,
        64'h626c7400_65707974,
        64'h2d756d6d_00617369,
        64'h2c766373_69720073,
        64'h75746174_73006765,
        64'h72006570_79745f65,
        64'h63697665_64007963,
        64'h6e657571_6572662d,
        64'h6b636f6c_63007963,
        64'h6e657571_6572662d,
        64'h65736162_656d6974,
        64'h00687461_702d7475,
        64'h6f647473_006c6564,
        64'h6f6d0065_6c626974,
        64'h61706d6f_6300736c,
        64'h6c65632d_657a6973,
        64'h2300736c_6c65632d,
        64'h73736572_64646123,
        64'h09000000_02000000,
        64'h02000000_02000000,
        64'h01000000_b5000000,
        64'h04000000_03000000,
        64'hffffffff_bf020000,
        64'h04000000_03000000,
        64'hffffffff_ae020000,
        64'h04000000_03000000,
        64'h01000000_a1020000,
        64'h04000000_03000000,
        64'h00000000_8a020000,
        64'h04000000_03000000,
        64'h08000000_79020000,
        64'h04000000_03000000,
        64'h08000000_69020000,
        64'h04000000_03000000,
        64'h00000000_55020000,
        64'h04000000_03000000,
        64'h00000000_43020000,
        64'h04000000_03000000,
        64'h00000000_31020000,
        64'h04000000_03000000,
        64'h00000000_21020000,
        64'h04000000_03000000,
        64'h00000100_00000000,
        64'h00000040_00000000,
        64'h67000000_10000000,
        64'h03000000_11020000,
        64'h00000000_03000000,
        64'h00000000_612e3030,
        64'h2e312d6f_6970672d,
        64'h7370782c_786e6c78,
        64'h1b000000_15000000,
        64'h03000000_02000000,
        64'h05020000_04000000,
        64'h03000000_00000030,
        64'h30303030_30303440,
        64'h6f697067_01000000,
        64'h02000000_00800000,
        64'h00000000_00000030,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h00007fe3_023e1800,
        64'hf3010000_06000000,
        64'h03000000_00000000,
        64'h03000000_52010000,
        64'h08000000_03000000,
        64'h03000000_41010000,
        64'h04000000_03000000,
        64'h006b726f_7774656e,
        64'h5b000000_08000000,
        64'h03000000_00687465,
        64'h2d637369_72776f6c,
        64'h1b000000_0c000000,
        64'h03000000_00000000,
        64'h30303030_30303033,
        64'h40687465_2d637369,
        64'h72776f6c_01000000,
        64'h02000000_02000000,
        64'he8010000_00000000,
        64'h03000000_e40c0000,
        64'he40c0000_d9010000,
        64'h08000000_03000000,
        64'h20bcbe00_c7010000,
        64'h04000000_03000000,
        64'h00000000_67000000,
        64'h04000000_03000000,
        64'h00000000_746f6c73,
        64'h2d697073_2d636d6d,
        64'h1b000000_0d000000,
        64'h03000000_00000030,
        64'h40636d6d_01000000,
        64'h04000000_b8010000,
        64'h04000000_03000000,
        64'h08000000_a1010000,
        64'h04000000_03000000,
        64'h01000000_90010000,
        64'h04000000_03000000,
        64'h01000000_80010000,
        64'h04000000_03000000,
        64'h00377865_746e696b,
        64'h74010000_08000000,
        64'h03000000_00100000,
        64'h00000000_00000020,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h02000000_02000000,
        64'h52010000_08000000,
        64'h03000000_03000000,
        64'h41010000_04000000,
        64'h03000000_00000000,
        64'h0f000000_04000000,
        64'h03000000_01000000,
        64'h00000000_04000000,
        64'h03000000_00612e30,
        64'h302e322d_6970732d,
        64'h7370782c_786e6c78,
        64'h00622e30_302e322d,
        64'h6970732d_7370782c,
        64'h786e6c78_1b000000,
        64'h28000000_03000000,
        64'h00000000_30303030,
        64'h30303032_40697073,
        64'h2d737078_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_0b010000,
        64'h08000000_03000000,
        64'h03000000_41010000,
        64'h04000000_03000000,
        64'h00100000_00000000,
        64'h00000018_00000000,
        64'h67000000_10000000,
        64'h03000000_07000000,
        64'h06000000_05000000,
        64'h04000000_52010000,
        64'h10000000_03000000,
        64'h00007265_6d69745f,
        64'h6270612c_706c7570,
        64'h1b000000_0f000000,
        64'h03000000_00003030,
        64'h30303030_38314072,
        64'h656d6974_01000000,
        64'h02000000_04000000,
        64'h67010000_04000000,
        64'h03000000_02000000,
        64'h5d010000_04000000,
        64'h03000000_01000000,
        64'h52010000_04000000,
        64'h03000000_03000000,
        64'h41010000_04000000,
        64'h03000000_00c20100,
        64'h33010000_04000000,
        64'h03000000_80f0fa02,
        64'h4b000000_04000000,
        64'h03000000_00100000,
        64'h00000000_00000010,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h00000000_61303535,
        64'h3631736e_1b000000,
        64'h09000000_03000000,
        64'h00000030_30303030,
        64'h30303140_74726175,
        64'h01000000_02000000,
        64'h03000000_b5000000,
        64'h04000000_03000000,
        64'h1e000000_28010000,
        64'h04000000_03000000,
        64'h07000000_15010000,
        64'h04000000_03000000,
        64'h00000004_00000000,
        64'h0000000c_00000000,
        64'h67000000_10000000,
        64'h03000000_09000000,
        64'h02000000_0b000000,
        64'h02000000_f7000000,
        64'h10000000_03000000,
        64'ha0000000_00000000,
        64'h03000000_00306369,
        64'h6c702c76_63736972,
        64'h1b000000_0c000000,
        64'h03000000_01000000,
        64'h8f000000_04000000,
        64'h03000000_00000000,
        64'h00000000_04000000,
        64'h03000000_00000000,
        64'h30303030_30306340,
        64'h72656c6c_6f72746e,
        64'h6f632d74_70757272,
        64'h65746e69_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_0b010000,
        64'h08000000_03000000,
        64'h00000c00_00000000,
        64'h00000002_00000000,
        64'h67000000_10000000,
        64'h03000000_07000000,
        64'h02000000_03000000,
        64'h02000000_f7000000,
        64'h10000000_03000000,
        64'h00000000_30746e69,
        64'h6c632c76_63736972,
        64'h1b000000_0d000000,
        64'h03000000_00000030,
        64'h30303030_30324074,
        64'h6e696c63_01000000,
        64'hf0000000_00000000,
        64'h03000000_00007375,
        64'h622d656c_706d6973,
        64'h00636f73_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h1f000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00636f73_01000000,
        64'h02000000_02000000,
        64'hd9000000_00000000,
        64'h03000000_00000074,
        64'h61656274_72616568,
        64'hc3000000_0a000000,
        64'h03000000_00000000,
        64'h01000000_01000000,
        64'hbd000000_0c000000,
        64'h03000000_00000064,
        64'h656c2d74_61656274,
        64'h72616568_01000000,
        64'h00000073_64656c2d,
        64'h6f697067_1b000000,
        64'h0a000000_03000000,
        64'h00000000_7364656c,
        64'h01000000_02000000,
        64'h00000040_00000000,
        64'h00000080_00000000,
        64'h67000000_10000000,
        64'h03000000_00007972,
        64'h6f6d656d_5b000000,
        64'h07000000_03000000,
        64'h00303030_30303030,
        64'h38407972_6f6d656d,
        64'h01000000_02000000,
        64'h02000000_02000000,
        64'h02000000_b5000000,
        64'h04000000_03000000,
        64'h00006374_6e692d75,
        64'h70632c76_63736972,
        64'h1b000000_0f000000,
        64'h03000000_a0000000,
        64'h00000000_03000000,
        64'h01000000_8f000000,
        64'h04000000_03000000,
        64'h00000000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h01000000_85000000,
        64'h00000000_03000000,
        64'h00003933_76732c76,
        64'h63736972_7c000000,
        64'h0b000000_03000000,
        64'h00006364_66616d69,
        64'h34367672_72000000,
        64'h0b000000_03000000,
        64'h00000076_63736972,
        64'h00656e61_69726120,
        64'h2c687465_1b000000,
        64'h12000000_03000000,
        64'h00000000_79616b6f,
        64'h6b000000_05000000,
        64'h03000000_00000000,
        64'h67000000_04000000,
        64'h03000000_00757063,
        64'h5b000000_04000000,
        64'h03000000_80f0fa02,
        64'h4b000000_04000000,
        64'h03000000_00000030,
        64'h40757063_01000000,
        64'h40787d01_38000000,
        64'h04000000_03000000,
        64'h00000000_0f000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00000000_73757063,
        64'h01000000_02000000,
        64'h00000030_30323531,
        64'h313a3030_30303030,
        64'h30314074_7261752f,
        64'h636f732f_2c000000,
        64'h1a000000_03000000,
        64'h00006e65_736f6863,
        64'h01000000_00657261,
        64'h622d656e_61697261,
        64'h2c687465_26000000,
        64'h10000000_03000000,
        64'h00766564_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h14000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00000000_01000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'he8080000_d2020000,
        64'h00000000_10000000,
        64'h11000000_28000000,
        64'h20090000_38000000,
        64'hf20b0000_edfe0dd0,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h46454443_42413938,
        64'h37363534_33323130,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h0000bdfd_c43e37fd,
        64'h10040413_47a29552,
        64'h414a8a33_b0003af3,
        64'h00f103a3_0ff7f793,
        64'h00044783_b0003a73,
        64'h94d2414a_8a33b000,
        64'h3af30154_0023b000,
        64'h3a73b701_c43e37fd,
        64'h10040413_47a29552,
        64'h414a8a33_b0003af3,
        64'h00f103a3_0ff7f793,
        64'h00044783_b0003a73,
        64'h94d2414a_8a33b000,
        64'h3af30154_0023b000,
        64'h3a73b709_c43e37fd,
        64'h10040413_47a29552,
        64'h414a8a33_b0003af3,
        64'h00f103a3_0ff7f793,
        64'h00044783_b0003a73,
        64'h94d2414a_8a33b000,
        64'h3af30154_0023b000,
        64'h3a73b569_00f102a3,
        64'h0ff7f793_37fd0051,
        64'h4783fc3e_838577e2,
        64'hb5450121_0323c781,
        64'h8ff97742_77e2b94d,
        64'hc63e2785_47b2b90f,
        64'hf0ef7502_b14ff0ef,
        64'h05050513_00001517,
        64'hba2ff0ef_6562b26f,
        64'hf0ef03a5_05130000,
        64'h1517f02a_ec260cf0,
        64'h44632781_47a24501,
        64'h4481c452_bc6ff0ef,
        64'h7502b4af_f0ef0365,
        64'h05130000_1517bd8f,
        64'hf0ef6562_b5cff0ef,
        64'h02050513_00001517,
        64'hf02aec26_0cf04363,
        64'h278147a2_45014481,
        64'hc44ebfcf_f0ef7502,
        64'hb80ff0ef_01c50513,
        64'h00001517_c0eff0ef,
        64'h6562b92f_f0ef0065,
        64'h05130000_1517f02a,
        64'hec260cf0_42632781,
        64'h47a24501_44819466,
        64'h90011402_c43e0640,
        64'h07934432_c3eff0ef,
        64'h7522bc2f_f0effe65,
        64'h05130000_1517c50f,
        64'hf0ef7502_bd4ff0ef,
        64'hfd850513_00001517,
        64'hc62ff0ef_6562be6f,
        64'hf0effd25_05130000,
        64'h1517cb6f_f0ef0ff5,
        64'h75136542_bfcff0ef,
        64'hfc850513_00001517,
        64'hcccff0ef_00514503,
        64'hc10ff0ef_fcc50513,
        64'h00001517_c1cff0ef,
        64'h07050513_00001517,
        64'he84ef462_f05a036a,
        64'h5c33416b_8b33b000,
        64'h3bf30124_89abb000,
        64'h3b734485_ec52414a,
        64'h8a33b000_3af31407,
        64'h86630ff7_f7930061,
        64'h4783b000_3a73fc62,
        64'hf84a0001_03230171,
        64'h02a3c6af_f0ef1fe5,
        64'h05130000_1517cf8f,
        64'hf0ef7522_c7cff0ef,
        64'h0a050513_00001517,
        64'hd0aff0ef_7502c8ef,
        64'hf0ef0925_05130000,
        64'h1517d1cf_f0ef6562,
        64'hca0ff0ef_08c50513,
        64'h00001517_d70ff0ef,
        64'h0ff57513_6542cb6f,
        64'hf0ef0825_05130000,
        64'h1517d86f_f0ef0041,
        64'h4503ccaf_f0ef0865,
        64'h05130000_1517cd6f,
        64'hf0ef1125_05130000,
        64'h1517e84e_f462f05a,
        64'h036a5c33_416b8b33,
        64'hb0003bf3_0124898b,
        64'hb0003b73_49019f84,
        64'h84930104_9493bfb4,
        64'h84930104_9493dfd4,
        64'h849bffff_04b7ec52,
        64'h414a8a33_b0003af3,
        64'hf7ed77c2_f83e83a1,
        64'h77c2fcf7_60e30ff7,
        64'hf7930041_470377c2,
        64'hbf31f83e_838577c2,
        64'h00f101a3_0ff7f793,
        64'h9fb98b85_00314703,
        64'h77c2b715_c43e37fd,
        64'h47a2bf19_c43e37fd,
        64'h47a2a82d_00f10223,
        64'h0ff7f793_77c2b000,
        64'h3a73f83e_5c47b783,
        64'h00001797_d7cff0ef,
        64'h31050513_00001517,
        64'he0aff0ef_7522d8ef,
        64'hf0ef1b25_05130000,
        64'h1517e1cf_f0ef7502,
        64'hda0ff0ef_1a450513,
        64'h00001517_e2eff0ef,
        64'h6562db2f_f0ef19e5,
        64'h05130000_1517e82f,
        64'hf0ef0ff5_75136542,
        64'hdc8ff0ef_19450513,
        64'h00001517_e98ff0ef,
        64'h00314503_ddcff0ef,
        64'h19850513_00001517,
        64'hde8ff0ef_18450513,
        64'h00001517_e84ef462,
        64'hf05a036a_5c33416b,
        64'h8b33b000_3bf30124,
        64'h89dbb000_3b7354fd,
        64'hec52414a_8a33b000,
        64'h3af3e7e9_77c2b000,
        64'h3a730001_01a3f85a,
        64'h0cf04963_278147a2,
        64'hc426f53f_f0ef4000,
        64'h05370ff0_05930ef0,
        64'h40632781_47a2c426,
        64'hf69ff0ef_0ff5f593,
        64'h40000537_65c26a0a,
        64'h0a137109_8993faa0,
        64'h0a9301f9_1c9303fb,
        64'h1c1303f0_0b93f9bf,
        64'hf0efb404_8493e76f,
        64'hf0ef6a61_69894905,
        64'h5b7d004c_54b720e5,
        64'h05130000_1517e4af,
        64'hf0efc602_e922e4e6,
        64'he8e2ecde_f0daf4d6,
        64'hf8d2fcce_e14ae526,
        64'hed060805_05130001,
        64'h03232005_859302fa,
        64'hf53765f1_000101a3,
        64'he83e0aa0_07937135,
        64'h808200e7_8623477d,
        64'h00078223_400007b7,
        64'h80820005_45038082,
        64'h00b50023_bbb9ee6f,
        64'hf0ef72a5_05130000,
        64'h1517bbc1_48450513,
        64'h00001517_f7eff0ef,
        64'h8526f02f_f0ef5865,
        64'h05130000_1517f0ef,
        64'hf0ef57a5_05130000,
        64'h1517bbe5_4ac50513,
        64'h00001517_fa6ff0ef,
        64'h8526f2af_f0ef5ae5,
        64'h05130000_1517f36f,
        64'hf0ef5a25_05130000,
        64'h1517c929_84aac3df,
        64'hf0ef9e0d_2605855a,
        64'h020aa583_028ab603,
        64'hf58ff0ef_78450513,
        64'h00001517_f3749de3,
        64'h08090913_08098993,
        64'hf70ff0ef_24855065,
        64'h05130000_1517ff49,
        64'h9be3847f_f0ef0a05,
        64'h000a4503_f8cff0ef,
        64'h7a850513_00001517,
        64'h81bff0ef_01093503,
        64'hfa0ff0ef_7ac50513,
        64'h00001517_82fff0ef,
        64'h00893503_fb4ff0ef,
        64'h7b050513_00001517,
        64'h843ff0ef_fb898a13,
        64'h00093503_fccff0ef,
        64'h7b850513_00001517,
        64'hff2a1be3_8a1ff0ef,
        64'h0a05000a_4503f909,
        64'h8a13feaf_f0ef7b65,
        64'h05130000_1517ff8a,
        64'h19e38bff_f0ef0a05,
        64'h0007c503_014c87b3,
        64'h4a0180bf_f0eff809,
        64'h8c937ba5_05130000,
        64'h15178dff_f0ef0ff4,
        64'hf513823f_f0ef7b65,
        64'h05130000_15174b91,
        64'h4c411005_1e630201,
        64'h09130801_099384aa,
        64'h8a8ad39f_f0ef850a,
        64'h46057101_04892583,
        64'h851ff0ef_5e450513,
        64'h00001517_89fff0ef,
        64'h4556863f_f0ef7d65,
        64'h05130000_15178b1f,
        64'hf0ef4546_875ff0ef,
        64'h7c850513_00001517,
        64'h903ff0ef_6526887f,
        64'hf0ef7ba5_05130000,
        64'h1517915f_f0ef7502,
        64'h899ff0ef_7bc50513,
        64'h00001517_927ff0ef,
        64'h65628abf_f0ef7b65,
        64'h05130000_15178f9f,
        64'hf0ef4552_8bdff0ef,
        64'h7b850513_00001517,
        64'h90bff0ef_45428cff,
        64'hf0ef7ba5_05130000,
        64'h151791df_f0ef4532,
        64'h8e1ff0ef_7bc50513,
        64'h00001517_92fff0ef,
        64'h45228f3f_f0ef7be5,
        64'h05130000_1517981f,
        64'hf0ef6502_905ff0ef,
        64'h7c050513_00001517,
        64'h911ff0ef_7ac50513,
        64'h00001517_bf5954f9,
        64'h921ff0ef_6b450513,
        64'h00001517_9afff0ef,
        64'h8526933f_f0ef7b65,
        64'h05130000_151793ff,
        64'hf0ef7aa5_05130000,
        64'h1517c905_84aa890a,
        64'he47ff0ef_850a4585,
        64'h46057101_95dff0ef,
        64'h7b050513_00001517,
        64'h80826125_6ca26c42,
        64'h6be27b02_7aa27a42,
        64'h79e26906_64a66446,
        64'h852660e6_fa040113,
        64'h54fd98bf_f0ef7b65,
        64'h05130000_1517c905,
        64'hdf3ff0ef_8b2a1080,
        64'he466e862_ec5ef456,
        64'hf852fc4e_e0cae4a6,
        64'hec86f05a_e8a2711d,
        64'hb7655479_80826169,
        64'h6baa6b4a_6aea7a0a,
        64'h79aa794a_74ea640e,
        64'h60ae8522_547d9d7f,
        64'hf0ef7da5_05130000,
        64'h1517c61f_f0efc65f,
        64'hf0efc69f_f0efc6df,
        64'hf0efc71f_f0efc75f,
        64'hf0efc79f_f0efc7df,
        64'hf0efa805_c83ff0ef,
        64'hc8dff0ef_45314581,
        64'h46054401_f93046e3,
        64'h20048493_19fda1ff,
        64'hf0ef8425_05130000,
        64'h2517e799_0369e7b3,
        64'h06891c63_90412901,
        64'h14428c49_cbbff0ef,
        64'h90410305_14130085,
        64'h151bcc9f_f0effc94,
        64'h1ae30404_0413ff7a,
        64'h17e3892a_f15ff0ef,
        64'h0a05854a_0007c583,
        64'h014407b3_04000b93,
        64'h4a01c6df_f0ef850a,
        64'h04000593_86224901,
        64'hff551ee3_d03ff0ef,
        64'he0048413_3e800b13,
        64'h0fe00a93_e9512004,
        64'h8493d1ff_f0ef4549,
        64'h85a20ff6_76130016,
        64'h66130015_161bf4df,
        64'hf0ef0ff4_7593f55f,
        64'hf0ef0ff5_f5930084,
        64'h559bf61f_f0ef0ff5,
        64'hf5930104_559bf6df,
        64'hf0ef4501_0184559b,
        64'hfee79be3_078500c6,
        64'h802300f1_06b30800,
        64'h0713567d_47810209,
        64'hd993842e_84aae55e,
        64'he95aed56_f152f94a,
        64'he586fd26_e1a20206,
        64'h1993f54e_71558082,
        64'h91411542_8d3d8ff9,
        64'h0057979b_17016709,
        64'h0107d79b_0105179b,
        64'h4105551b_0105151b,
        64'h8d2d00c5_95138da9,
        64'h893d0045_d51b8da9,
        64'h91411542_8d5d0522,
        64'h0085579b_808207f5,
        64'h75138d2d_00451593,
        64'h8d2d8d3d_0045d51b,
        64'h0075d79b_8de98082,
        64'h0141853e_640260a2,
        64'h57f5e111_4781f89f,
        64'hf0efc511_57f9efbf,
        64'hf0efc911_57fdeb7f,
        64'hf0effc6d_e0bff0ef,
        64'h347d4429_b95ff0ef,
        64'h98050513_00002517,
        64'hc8fff0ef_e022e406,
        64'h11418082_61050015,
        64'h351364a2_644260e2,
        64'h0004051b_fc940ce3,
        64'he3fff0ef_eb5ff0ef,
        64'h9a850513_00002517,
        64'h85aa842a_e59ff0ef,
        64'h02900513_400005b7,
        64'h07700613_fbdff0ef,
        64'h4485e822_ec06e426,
        64'h11018082_01410015,
        64'h3513157d_640260a2,
        64'h0004051b_ef5ff0ef,
        64'h9e250513_85a20000,
        64'h2517e91f_f0ef842a,
        64'he9dff0ef_e022e406,
        64'h03700513_45810650,
        64'h06131141_80826105,
        64'h690264a2_644260e2,
        64'h00153513_f5650513,
        64'h0004051b_01249863,
        64'h88bd00f9_1b634501,
        64'h4785ed1f_f0efed5f,
        64'hf0ef842a_edbff0ef,
        64'h84aaee1f_f0efee5f,
        64'hf0efee9f_f0ef892a,
        64'hef5ff0ef_e04ae426,
        64'he822ec06_45211aa0,
        64'h05930870_06131101,
        64'hbfcd4501_80826105,
        64'h690264a2_644260e2,
        64'h4505f8bf_f0ef4585,
        64'ha7050513_00002517,
        64'hfe9915e3_c00df2df,
        64'hf0ef892a_347df3bf,
        64'hf0ef4501_45810950,
        64'h06134485_71040413,
        64'he04aec06_e4266409,
        64'he8221101_b9c96105,
        64'ha6850513_00002517,
        64'h60e26442_da9ff0ef,
        64'h852e65a2_cedff0ef,
        64'hab050513_00002517,
        64'hcf9ff0ef_8522cfff,
        64'hf0efe42e_ec06ab65,
        64'h05130000_2517842a,
        64'he8221101_80826145,
        64'h64e27402_70a2f47d,
        64'h147d0007_d4634187,
        64'hd79b0185_179bfadf,
        64'hf0efeb7f_f0ef8532,
        64'h06400413_6622ec3f,
        64'hf0ef0ff4_7513ecbf,
        64'hf0ef0ff5_75130084,
        64'h551bed7f_f0ef0ff5,
        64'h75130104_551bee3f,
        64'hf0ef0184_551beebf,
        64'hf0ef0404_e513fedf,
        64'hf0ef84aa_842eec26,
        64'hf022e432_f4067179,
        64'hb7090ff0_05138082,
        64'h557db7d9_00d70023,
        64'h078500f6_073306c8,
        64'h2683ff69_8b055178,
        64'hb77dd6b8_07850007,
        64'h470300f5_07338082,
        64'h4501d3b8_4719dbb8,
        64'h577d2000_07b702b6,
        64'he1630007_869b2000,
        64'h08372000_0537fff5,
        64'h8b85537c_20000737,
        64'hd3b82000_07b71060,
        64'h0713fff5_37fd0001,
        64'h03200793_04b76163,
        64'h0007871b_47812000,
        64'h06b7dbb8_57792000,
        64'h07b706b7_ee631000,
        64'h07938082_610564a2,
        64'hd3b84719_dbb86442,
        64'h60e20ff4_7513577d,
        64'h200007b7_e25ff0ef,
        64'hbb850513_00002517,
        64'heb3ff0ef_91011502,
        64'h4088e3bf_f0efbd65,
        64'h05130000_2517e395,
        64'h8b852401_53fc57e0,
        64'hff658b05_06478493,
        64'h53f8d3b8_10600713,
        64'h200007b7_fff537fd,
        64'h00010640_0793d7a8,
        64'hdbb85779_e426e822,
        64'hec062000_07b71101,
        64'hbdbd6105_c0450513,
        64'h00002517_64a260e2,
        64'h6442d03c_4799e97f,
        64'hf0efc2a5_05130000,
        64'h2517f25f_f0ef9101,
        64'h02049513_2481eaff,
        64'hf0efc225_05130000,
        64'h25175064_d03c1660,
        64'h0793ec3f_f0efc565,
        64'h05130000_2517f51f,
        64'hf0ef9101_02049513,
        64'h2481edbf_f0efc4e5,
        64'h05130000_25175064,
        64'hd03c1040_07932000,
        64'h0437fff5_37fd0001,
        64'h47a9c3b8_47292000,
        64'h07b7f03f_f0efe426,
        64'he822ec06_c6e50513,
        64'h11010000_25178082,
        64'h25014108_8082c10c,
        64'h80826105_60e2ecff,
        64'hf0ef0091_4503ed7f,
        64'hf0ef0081_4503f55f,
        64'hf0efec06_002c1101,
        64'h80826145_694264e2,
        64'h740270a2_fe9410e3,
        64'hef9ff0ef_00914503,
        64'hf01ff0ef_34610081,
        64'h4503f81f_f0ef0ff5,
        64'h7513002c_00895533,
        64'h54e10380_0413892a,
        64'hf406e84a_ec26f022,
        64'h71798082_61456942,
        64'h64e27402_70a2fe94,
        64'h10e3f3bf_f0ef0091,
        64'h4503f43f_f0ef3461,
        64'h00814503_fc3ff0ef,
        64'h0ff57513_002c0089,
        64'h553b54e1_4461892a,
        64'hf406e84a_ec26f022,
        64'h71798082_00f58023,
        64'h0007c783_00e580a3,
        64'h97aa8111_00074703,
        64'h973e00f5_7713e6e7,
        64'h87930000_1797b7f5,
        64'h0405f93f_f0ef8082,
        64'h01416402_60a2e509,
        64'h00044503_842ae406,
        64'he0221141_808200e7,
        64'h88230200_071300e7,
        64'h8423fc70_071300e7,
        64'h8623470d_00a78223,
        64'h0ff57513_00e78023,
        64'h0085551b_0ff57713,
        64'h00e78623_f8000713,
        64'h00078223_100007b7,
        64'h02b5553b_0045959b,
        64'h808200a7_0023dfe5,
        64'h0207f793_01474783,
        64'h10000737_80820205,
        64'h75130147_c5031000,
        64'h07b78082_00054503,
        64'h808200b5_00238082,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00048067_01f49493,
        64'h0010049b_08458593,
        64'h00001597_f1402573,
        64'hff24c6e3_4009091b,
        64'h02000937_00448493,
        64'hfe091ee3_0004a903,
        64'h00092023_00990933,
        64'h00291913_f1402973,
        64'h020004b7_fe090ae3,
        64'h00897913_34402973,
        64'h10500073_ff24c6e3,
        64'h4009091b_02000937,
        64'h00448493_0124a023,
        64'h00100913_020004b7,
        64'h295000ef_01a11113,
        64'h0210011b_03249663,
        64'hf1402973_00000493,
        64'h30491073_00800913
    };

    logic [$clog2(RomSize)-1:0] addr_q;

    always_ff @(posedge clk_i) begin
        if (req_i) begin
            addr_q <= addr_i[$clog2(RomSize)-1+3:3];
        end
    end

    // this prevents spurious Xes from propagating into
    // the speculative fetch stage of the core
    assign rdata_o = (addr_q < RomSize) ? mem[addr_q] : '0;
endmodule
